netcdf ulong_3d {
dimensions:
	dim_0 = 2 ;
	dim_1 = 10 ;
	dim_2 = 5 ;
variables:
	int values(dim_0, dim_1, dim_2) ;
		values:valid_min = -2147483648 ;
		values:valid_max = 2147483647 ;
data:

 values =
  -2147483648, _, -2147483646, -2147483645, -2147483644,
  _, -2147483646, -2147483645, -2147483644, -2147483643,
  -2147483646, -2147483645, -2147483644, -2147483643, -2147483642,
  -2147483645, -2147483644, -2147483643, -2147483642, -2147483641,
  -2147483644, -2147483643, -2147483642, -2147483641, -2147483640,
  -2147483643, -2147483642, -2147483641, -2147483640, -2147483639,
  -2147483642, -2147483641, -2147483640, -2147483639, -2147483638,
  -2147483641, -2147483640, -2147483639, -2147483638, -2147483637,
  -2147483640, -2147483639, -2147483638, -2147483637, -2147483636,
  -2147483639, -2147483638, -2147483637, -2147483636, -2147483635,
  _, -2147483646, -2147483645, -2147483644, -2147483643,
  -2147483646, -2147483645, -2147483644, -2147483643, -2147483642,
  -2147483645, -2147483644, -2147483643, -2147483642, -2147483641,
  -2147483644, -2147483643, -2147483642, -2147483641, -2147483640,
  -2147483643, -2147483642, -2147483641, -2147483640, -2147483639,
  -2147483642, -2147483641, -2147483640, -2147483639, -2147483638,
  -2147483641, -2147483640, -2147483639, -2147483638, -2147483637,
  -2147483640, -2147483639, -2147483638, -2147483637, -2147483636,
  -2147483639, -2147483638, -2147483637, -2147483636, -2147483635,
  -2147483638, -2147483637, -2147483636, -2147483635, -2147483634 ;
}
