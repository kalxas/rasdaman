netcdf double_4d_transpose_import {
dimensions:
	dim_0 = 2 ;
	dim_1 = 2 ;
	dim_2 = 5 ;
	dim_3 = 10 ;
variables:
	double values(dim_0, dim_1, dim_2, dim_3) ;
		values:missing_value = "NaN" ;
data:

 values =
  1, 6, 11, 16, 21, 26, 31, 36, 41, 46,
  2, 7, 12, 17, 22, 27, 32, 37, 42, 47,
  3, 8, 13, 18, 23, 28, 33, 38, 43, 48,
  4, 9, 14, 19, 24, 29, 34, 39, 44, 49,
  5, 10, 15, 20, 25, 30, 35, 40, 45, 50,
  51, 56, 61, 66, 71, 76, 81, 86, 91, 96,
  52, 57, 62, 67, 72, 77, 82, 87, 92, 97,
  53, 58, 63, 68, 73, 78, 83, 88, 93, 98,
  54, 59, 64, 69, 74, 79, 84, 89, 94, 99,
  55, 60, 65, 70, 75, 80, 85, 90, 95, 100,
  101, 106, 111, 116, 121, 126, 131, 136, 141, 146,
  102, 107, 112, 117, 122, 127, 132, 137, 142, 147,
  103, 108, 113, 118, 123, 128, 133, 138, 143, 148,
  104, 109, 114, 119, 124, 129, 134, 139, 144, 149,
  105, 110, 115, 120, 125, 130, 135, 140, 145, 150,
  151, 156, 161, 166, 171, 176, 181, 186, 191, 196,
  152, 157, 162, 167, 172, 177, 182, 187, 192, 197,
  153, 158, 163, 168, 173, 178, 183, 188, 193, 198,
  154, 159, 164, 169, 174, 179, 184, 189, 194, 199,
  155, 160, 165, 170, 175, 180, 185, 190, 195, 200 ;
}
