netcdf long_3d {
dimensions:
	dim_0 = 3 ;
	dim_1 = 10 ;
	dim_2 = 5 ;
variables:
	int values(dim_0, dim_1, dim_2) ;
		values:valid_min = -2147483648 ;
		values:valid_max = 2147483647 ;
data:

 values =
  1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15,
  16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30,
  31, 32, 33, 34, 35,
  36, 37, 38, 39, 40,
  41, 42, 43, 44, 45,
  46, 47, 48, 49, 50,
  51, 52, 53, 54, 55,
  56, 57, 58, 59, 60,
  61, 62, 63, 64, 65,
  66, 67, 68, 69, 70,
  71, 72, 73, 74, 75,
  76, 77, 78, 79, 80,
  81, 82, 83, 84, 85,
  86, 87, 88, 89, 90,
  91, 92, 93, 94, 95,
  96, 97, 98, 99, 100,
  101, 102, 103, 104, 105,
  106, 107, 108, 109, 110,
  111, 112, 113, 114, 115,
  116, 117, 118, 119, 120,
  121, 122, 123, 124, 125,
  126, 127, 128, 129, 130,
  131, 132, 133, 134, 135,
  136, 137, 138, 139, 140,
  141, 142, 143, 144, 145,
  146, 147, 148, 149, 150 ;
}
