netcdf ushort_4d {
dimensions:
	dim_0 = 2 ;
	dim_1 = 2 ;
	dim_2 = 10 ;
	dim_3 = 5 ;
variables:
	int values(dim_0, dim_1, dim_2, dim_3) ;
		values:valid_min = 0 ;
		values:valid_max = 65535 ;
data:

 values =
  32768, 32769, 32770, 32771, 32772,
  32769, 32770, 32771, 32772, 32773,
  32770, 32771, 32772, 32773, 32774,
  32771, 32772, 32773, 32774, 32775,
  32772, 32773, 32774, 32775, 32776,
  32773, 32774, 32775, 32776, 32777,
  32774, 32775, 32776, 32777, 32778,
  32775, 32776, 32777, 32778, 32779,
  32776, 32777, 32778, 32779, 32780,
  32777, 32778, 32779, 32780, 32781,
  32769, 32770, 32771, 32772, 32773,
  32770, 32771, 32772, 32773, 32774,
  32771, 32772, 32773, 32774, 32775,
  32772, 32773, 32774, 32775, 32776,
  32773, 32774, 32775, 32776, 32777,
  32774, 32775, 32776, 32777, 32778,
  32775, 32776, 32777, 32778, 32779,
  32776, 32777, 32778, 32779, 32780,
  32777, 32778, 32779, 32780, 32781,
  32778, 32779, 32780, 32781, 32782,
  32769, 32770, 32771, 32772, 32773,
  32770, 32771, 32772, 32773, 32774,
  32771, 32772, 32773, 32774, 32775,
  32772, 32773, 32774, 32775, 32776,
  32773, 32774, 32775, 32776, 32777,
  32774, 32775, 32776, 32777, 32778,
  32775, 32776, 32777, 32778, 32779,
  32776, 32777, 32778, 32779, 32780,
  32777, 32778, 32779, 32780, 32781,
  32778, 32779, 32780, 32781, 32782,
  32770, 32771, 32772, 32773, 32774,
  32771, 32772, 32773, 32774, 32775,
  32772, 32773, 32774, 32775, 32776,
  32773, 32774, 32775, 32776, 32777,
  32774, 32775, 32776, 32777, 32778,
  32775, 32776, 32777, 32778, 32779,
  32776, 32777, 32778, 32779, 32780,
  32777, 32778, 32779, 32780, 32781,
  32778, 32779, 32780, 32781, 32782,
  32779, 32780, 32781, 32782, 32783 ;
}
