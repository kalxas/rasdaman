netcdf octet_4d_transpose_import {
dimensions:
	dim_0 = 1 ;
	dim_1 = 2 ;
	dim_2 = 5 ;
	dim_3 = 10 ;
variables:
	byte values(dim_0, dim_1, dim_2, dim_3) ;
		values:valid_min = -128b ;
		values:valid_max = 127b ;
data:

 values =
  -1, 6, 11, 16, 21, 26, 31, 36, 41, 46,
  2, 7, 12, 17, 22, 27, 32, 37, 42, 47,
  3, 8, 13, 18, 23, 28, 33, 38, 43, 48,
  4, 9, 14, 19, 24, 29, 34, 39, 44, 49,
  5, 10, 15, 20, 25, 30, 35, 40, 45, 50,
  51, 56, 61, 66, 71, 76, 81, 86, 91, 96,
  52, 57, 62, 67, 72, 77, 82, 87, 92, 97,
  53, 58, 63, 68, 73, 78, 83, 88, 93, 98,
  54, 59, 64, 69, 74, 79, 84, 89, 94, 99,
  55, 60, 65, 70, 75, 80, 85, 90, 95, 100 ;
}
