netcdf char_3d {
dimensions:
	dim_0 = 2 ;
	dim_1 = 10 ;
	dim_2 = 5 ;
variables:
	short values(dim_0, dim_1, dim_2) ;
		values:valid_min = 0s ;
		values:valid_max = 255s ;
data:

 values =
  128, 129, 130, 131, 132,
  129, 130, 131, 132, 133,
  130, 131, 132, 133, 134,
  131, 132, 133, 134, 135,
  132, 133, 134, 135, 136,
  133, 134, 135, 136, 137,
  134, 135, 136, 137, 138,
  135, 136, 137, 138, 139,
  136, 137, 138, 139, 140,
  137, 138, 139, 140, 141,
  129, 130, 131, 132, 133,
  130, 131, 132, 133, 134,
  131, 132, 133, 134, 135,
  132, 133, 134, 135, 136,
  133, 134, 135, 136, 137,
  134, 135, 136, 137, 138,
  135, 136, 137, 138, 139,
  136, 137, 138, 139, 140,
  137, 138, 139, 140, 141,
  138, 139, 140, 141, 142 ;
}
