netcdf octet_3d_json_export {
dimensions:
	time = 2 ;
	lat = 10 ;
	lon = 5 ;
variables:
	byte tos(time, lat, lon) ;
		tos:valid_min = -128b ;
		tos:valid_max = 127b ;
		tos:cell_methods = "time: mean (interval: 30 minutes)" ;
		tos:history = " At 16:37:23 on 01/11/2005: CMOR altered the data in the following ways: added 2.73150E+02 to yield output units; Cyclical dimension was output starting at a different lon;" ;
		tos:long_name = "Sea Surface Temperature" ;
		tos:missing_value = 1.e+20 ;
		tos:original_name = "sosstsst" ;
		tos:original_units = "degC" ;
		tos:standard_name = "sea_surface_temperature" ;
		tos:units = "K" ;
	double lat(lat) ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
		lat:long_name = "latitude" ;
		lat:original_units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(lon) ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
		lon:long_name = "longitude" ;
		lon:original_units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:calendar = "360_day" ;
		time:long_name = "time" ;
		time:original_units = "seconds since 2001-1-1" ;
		time:standard_name = "time" ;
		time:units = "days since 2001-1-1" ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:cmor_version = 0.96 ;
		:comment = "Test drive" ;
		:contact = "Sebastien Denvil, sebastien.denvil@ipsl.jussieu.fr" ;
		:experiment_id = "SRES A2 experiment" ;
		:history = "YYYY/MM/JJ: data generated; YYYY/MM/JJ+1 data transformed At 16:37:23 on 01/11/2005, CMOR rewrote data to comply with CF standards and IPCC Fourth Assessment requirements" ;
		:institution = "IPSL (Institut Pierre Simon Laplace, Paris, France)" ;
		:project_id = "IPCC Fourth Assessment" ;
		:realization = 1LL ;
		:references = "Dufresne et al, Journal of Climate, 2015, vol XX, p 136" ;
		:source = "IPSL-CM4_v1 (2003) : atmosphere : LMDZ (IPSL-CM4_IPCC, 96x71x19), ocean ORCA2 (ipsl_cm4_v1_8, 2x2L31); sea ice LIM (ipsl_cm4_v" ;
		:table_id = "Table O1 (13 November 2004)" ;
		:title = "IPSL model output prepared for IPCC Fourth Assessment SRES A2 experiment" ;
data:

 tos =
  -1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15,
  16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30,
  31, 32, 33, 34, 35,
  36, 37, 38, 39, 40,
  41, 42, 43, 44, 45,
  46, 47, 48, 49, 50,
  51, 52, 53, 54, 55,
  56, 57, 58, 59, 60,
  61, 62, 63, 64, 65,
  66, 67, 68, 69, 70,
  71, 72, 73, 74, 75,
  76, 77, 78, 79, 80,
  81, 82, 83, 84, 85,
  86, 87, 88, 89, 90,
  91, 92, 93, 94, 95,
  96, 97, 98, 99, 100 ;

 lat = -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, -70.5 ;

 lon = 1, 3, 5, 7, 9 ;

 time = 15, 45 ;
}
