netcdf octet_3d_json_import_subsetDomain {
dimensions:
	dim_0 = 1 ;
	dim_1 = 10 ;
	dim_2 = 3 ;
variables:
	byte values(dim_0, dim_1, dim_2) ;
		values:valid_min = -128b ;
		values:valid_max = 127b ;
data:

 values =
  -1, 2, 3,
  6, 7, 8,
  11, 12, 13,
  16, 17, 18,
  21, 22, 23,
  26, 27, 28,
  31, 32, 33,
  36, 37, 38,
  41, 42, 43,
  46, 47, 48 ;
}
