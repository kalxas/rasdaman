netcdf ulong_3d {
dimensions:
	dim_0 = 2 ;
	dim_1 = 10 ;
	dim_2 = 5 ;
variables:
	uint values(dim_0, dim_1, dim_2) ;
		values:valid_min = 0U ;
		values:valid_max = 4294967295U ;
data:

 values =
  2147483648, 2147483649, 2147483650, 2147483651, 2147483652,
  2147483649, 2147483650, 2147483651, 2147483652, 2147483653,
  2147483650, 2147483651, 2147483652, 2147483653, 2147483654,
  2147483651, 2147483652, 2147483653, 2147483654, 2147483655,
  2147483652, 2147483653, 2147483654, 2147483655, 2147483656,
  2147483653, 2147483654, 2147483655, 2147483656, 2147483657,
  2147483654, 2147483655, 2147483656, 2147483657, 2147483658,
  2147483655, 2147483656, 2147483657, 2147483658, 2147483659,
  2147483656, 2147483657, 2147483658, 2147483659, 2147483660,
  2147483657, 2147483658, 2147483659, 2147483660, 2147483661,
  2147483649, 2147483650, 2147483651, 2147483652, 2147483653,
  2147483650, 2147483651, 2147483652, 2147483653, 2147483654,
  2147483651, 2147483652, 2147483653, 2147483654, 2147483655,
  2147483652, 2147483653, 2147483654, 2147483655, 2147483656,
  2147483653, 2147483654, 2147483655, 2147483656, 2147483657,
  2147483654, 2147483655, 2147483656, 2147483657, 2147483658,
  2147483655, 2147483656, 2147483657, 2147483658, 2147483659,
  2147483656, 2147483657, 2147483658, 2147483659, 2147483660,
  2147483657, 2147483658, 2147483659, 2147483660, 2147483661,
  2147483658, 2147483659, 2147483660, 2147483661, 2147483662 ;
}
