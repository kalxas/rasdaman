netcdf float_3d {
dimensions:
	dim_0 = 3 ;
	dim_1 = 10 ;
	dim_2 = 5 ;
variables:
	float values(dim_0, dim_1, dim_2) ;
		values:missing_value = "NaNf" ;
data:

 values =
  1.5, 2.5, 3.5, 4.5, 5.5,
  6.5, 7.5, 8.5, 9.5, 10.5,
  11.5, 12.5, 13.5, 14.5, 15.5,
  16.5, 17.5, 18.5, 19.5, 20.5,
  21.5, 22.5, 23.5, 24.5, 25.5,
  26.5, 27.5, 28.5, 29.5, 30.5,
  31.5, 32.5, 33.5, 34.5, 35.5,
  36.5, 37.5, 38.5, 39.5, 40.5,
  41.5, 42.5, 43.5, 44.5, 45.5,
  46.5, 47.5, 48.5, 49.5, 50.5,
  51.5, 52.5, 53.5, 54.5, 55.5,
  56.5, 57.5, 58.5, 59.5, 60.5,
  61.5, 62.5, 63.5, 64.5, 65.5,
  66.5, 67.5, 68.5, 69.5, 70.5,
  71.5, 72.5, 73.5, 74.5, 75.5,
  76.5, 77.5, 78.5, 79.5, 80.5,
  81.5, 82.5, 83.5, 84.5, 85.5,
  86.5, 87.5, 88.5, 89.5, 90.5,
  91.5, 92.5, 93.5, 94.5, 95.5,
  96.5, 97.5, 98.5, 99.5, 100.5,
  101.5, 102.5, 103.5, 104.5, 105.5,
  106.5, 107.5, 108.5, 109.5, 110.5,
  111.5, 112.5, 113.5, 114.5, 115.5,
  116.5, 117.5, 118.5, 119.5, 120.5,
  121.5, 122.5, 123.5, 124.5, 125.5,
  126.5, 127.5, 128.5, 129.5, 130.5,
  131.5, 132.5, 133.5, 134.5, 135.5,
  136.5, 137.5, 138.5, 139.5, 140.5,
  141.5, 142.5, 143.5, 144.5, 145.5,
  146.5, 147.5, 148.5, 149.5, 150.5 ;
}
